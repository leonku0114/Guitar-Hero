module HexDriver (input  [6:0]  In0,
                  output logic [13:0]  Out0);
	
	always_comb
	begin
//		unique case (In0)
//	 	   4'b0000   : Out0 = 7'b1000000; // '0'
//	 	   4'b0001   : Out0 = 7'b1111001; // '1'
//		   4'b0010   : Out0 = 7'b0100100; // '2'
//	 	   4'b0011   : Out0 = 7'b0110000; // '3'
//	 	   4'b0100   : Out0 = 7'b0011001; // '4'
//		   4'b0101   : Out0 = 7'b0010010; // '5'
//	 	   4'b0110   : Out0 = 7'b0000010; // '6'
//	 	   4'b0111   : Out0 = 7'b1111000; // '7'
//	 	   4'b1000   : Out0 = 7'b0000000; // '8'
//		   4'b1001   : Out0 = 7'b0010000; // '9'
//	 	   4'b1010   : Out0 = 7'b0001000; // 'A'
//	 	   4'b1011   : Out0 = 7'b0000011; // 'b'
//	 	   4'b1100   : Out0 = 7'b1000110; // 'C'
//		   4'b1101   : Out0 = 7'b0100001; // 'd'
//	 	   4'b1110   : Out0 = 7'b0000110; // 'E'
//	 	   4'b1111   : Out0 = 7'b0001110; // 'F'
//	 	   default   : Out0 = 7'bX;
//	  	 endcase


unique case (In0)
	 	   7'b0000000   : Out0 = 14'b00000001110111; // '0'
	 	   7'b0000001   : Out0 = 14'b00000000010010; // '1'
		   7'b0000010   : Out0 = 14'b00000001011101; // '2'
	 	   7'b0000011   : Out0 = 14'b00000001011011; // '3'
	 	   7'b0000100   : Out0 = 14'b00000000111010; // '4'
		   7'b0000101   : Out0 = 14'b00000001101011; // '5'
	 	   7'b0000110   : Out0 = 14'b00000001101111; // '6'
	 	   7'b0000111   : Out0 = 14'b00000001010010; // '7'
	 	   7'b0001000   : Out0 = 14'b00000001111111; // '8'
		   7'b0001001   : Out0 = 14'b00000001111010; // '9'
			
	 	   7'b0001010   : Out0 = 14'b00100101110111; // '10'
	 	   7'b0001011   : Out0 = 14'b00100100010010; // '11'
	 	   7'b0001100   : Out0 = 14'b00100101011101; // '12'
		   7'b0001101   : Out0 = 14'b00100101011011; // '13'
	 	   7'b0001110   : Out0 = 14'b00100100111010; // '14'
	 	   7'b0001111   : Out0 = 14'b00100101101011; // '15'
			7'b0010000   : Out0 = 14'b00100101101111; // '16'
			7'b0010001   : Out0 = 14'b00100101010010; // '17'
			7'b0010010   : Out0 = 14'b00100101111111; // '18'
			7'b0010011   : Out0 = 14'b00100101111010; // '19'
			
			7'b0010100   : Out0 = 14'b10111011110111; // '20'0010100
			7'b0010101   : Out0 = 14'b10111010010010; // '21'
			7'b0010110   : Out0 = 14'b10111011011101; // '22'
			7'b0010111   : Out0 = 14'b10111011011011; // '23'
			7'b0011000   : Out0 = 14'b10111010111010; // '24'
			7'b0011001   : Out0 = 14'b10111011101011; // '25'
			7'b0011010   : Out0 = 14'b10111011101111; // '26'
			7'b0011011   : Out0 = 14'b10111011010010; // '27'
			7'b0011100   : Out0 = 14'b10111011111111; // '28'
			7'b0011101   : Out0 = 14'b10111011111010; // '29'
			
			7'b0011110   : Out0 = 14'b10110111110111; // '30'
			7'b0011111   : Out0 = 14'b10110110010010; // '31'			
			7'b0100000   : Out0 = 14'b10110111011101; // '32'
			7'b0100001   : Out0 = 14'b10110111011011; // '33'
			7'b0100010   : Out0 = 14'b10110110111010; // '34'
			7'b0100011   : Out0 = 14'b10110111101011; // '35'
			7'b0100100   : Out0 = 14'b10110111101111; // '36'
			7'b0100101   : Out0 = 14'b10110111010010; // '37'
			7'b0100110   : Out0 = 14'b10110111111111; // '38'
			7'b0100111   : Out0 = 14'b10110111111010; // '39'
			
			
			7'b0101000   : Out0 = 14'b01110101110111; // '40'
			7'b0101001   : Out0 = 14'b01110100010010; // '41'			
			7'b0101010   : Out0 = 14'b01110101011101; // '42'
			7'b0101011   : Out0 = 14'b01110101011011; // '43'
			7'b0101100   : Out0 = 14'b01110100111010; // '44'
			7'b0101101   : Out0 = 14'b01110101101011; // '45'
			7'b0101110   : Out0 = 14'b01110101101111; // '46'
			7'b0101111   : Out0 = 14'b01110101010010; // '47'
			7'b0110000   : Out0 = 14'b01110101111111; // '48'
			7'b0110001   : Out0 = 14'b01110101111010; // '49'
			
			7'b0110010   : Out0 = 14'b11010111110111; // '50'
			7'b0110011   : Out0 = 14'b11010110010010; // '51'			
			7'b0110100   : Out0 = 14'b11010111011101; // '52'
			7'b0110101   : Out0 = 14'b11010111011011; // '53'
			7'b0110110   : Out0 = 14'b11010110111010; // '54'
			7'b0110111   : Out0 = 14'b11010111101011; // '55'
			7'b0111000   : Out0 = 14'b11010111101111; // '56'
			7'b0111001   : Out0 = 14'b11010111010010; // '57'
			7'b0111010   : Out0 = 14'b11010111111111; // '58'
			7'b0111011   : Out0 = 14'b11010111111010; // '59'
			
			7'b0111100   : Out0 = 14'b11011111110111; // '60'
			7'b0111101   : Out0 = 14'b11011110010010; // '61'			
			7'b0111110   : Out0 = 14'b11011111011101; // '62'
			7'b0111111   : Out0 = 14'b11011111011011; // '63'
			7'b1000000   : Out0 = 14'b11011110111010; // '64'
			7'b1000001   : Out0 = 14'b11011111101011; // '65'
			7'b1000010   : Out0 = 14'b11011111101111; // '66'
			7'b1000011   : Out0 = 14'b11011111010010; // '67'
			7'b1000100   : Out0 = 14'b11011111111111; // '68'
			7'b1000101   : Out0 = 14'b11011111111010; // '69'
			
			7'b1000110   : Out0 = 14'b10100101110111; // '70'
			7'b1000111   : Out0 = 14'b10100100010010; // '71'			
			7'b1001000   : Out0 = 14'b10100101011101; // '72'
			7'b1001001   : Out0 = 14'b10100101011011; // '73'
			7'b1001010   : Out0 = 14'b10100100111010; // '74'
			7'b1001011   : Out0 = 14'b10100101101011; // '75'
			7'b1001100   : Out0 = 14'b10100101101111; // '76'
			7'b1001101   : Out0 = 14'b10100101010010; // '77'
			7'b1001110   : Out0 = 14'b10100101111111; // '78'
			7'b1001111   : Out0 = 14'b10100101111010; // '79'
			
			7'b1010000   : Out0 = 14'b11111111110111; // '80'
			7'b1010001   : Out0 = 14'b11111110010010; // '81'			
			7'b1010010   : Out0 = 14'b11111111011101; // '82'
			7'b1010011   : Out0 = 14'b11111111011011; // '83'
			7'b1010100   : Out0 = 14'b11111110111010; // '84'
			7'b1010101   : Out0 = 14'b11111111101011; // '85'
			7'b1010110   : Out0 = 14'b11111111101111; // '86'
			7'b1010111   : Out0 = 14'b11111111010010; // '87'
			7'b1011000   : Out0 = 14'b11111110010010; // '88'
			7'b1011001   : Out0 = 14'b11111111111010; // '89'
	 	   default   : Out0 = 7'bX;
	  	 endcase
	end

endmodule